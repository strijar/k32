--
--  Copyright 2015-2026 Oleg Belousov <belousov.oleg@gmail.com>,
--
--  All rights reserved.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--    1. Redistributions of source code must retain the above copyright notice,
--       this list of conditions and the following disclaimer.
-- 
--    2. Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.k32_pkg.all;

entity ram is
    generic (
	addr_bits	: integer := 5;
	data_bits	: integer := 16
    );
    port (
	clk	: in std_logic;
	rst	: in std_logic;

	a_addr	: in std_logic_vector(addr_bits-1 downto 0);
	a_din	: in std_logic_vector(data_bits-1 downto 0);
	a_dout	: out std_logic_vector(data_bits-1 downto 0);
        a_we	: in std_logic;

	b_en	: in std_logic;
	b_addr	: in std_logic_vector(addr_bits-1 downto 0);
	b_din	: in std_logic_vector(data_bits-1 downto 0);
	b_dout	: out std_logic_vector(data_bits-1 downto 0);
        b_we	: in std_logic_vector(3 downto 0)
    );
end ram;

architecture rtl of ram is

type ram_type is array(natural range 0 to (2**(addr_bits))-1) of std_logic_vector(data_bits-1 downto 0);

signal a_addr_word	: std_logic_vector(addr_bits-1 downto 2) := (others => '0');
signal b_addr_word	: std_logic_vector(addr_bits-1 downto 2) := (others => '0');

signal ram : ram_type :=
(
0000 => x"000003A0",	--0000
0001 => x"000009E8",	--0004

0008 => x"00000000",	--0020
0009 => x"00000000",	--0024
0010 => x"00000000",	--0028
0011 => x"00000000",	--002C
0012 => x"00000000",	--0030
0013 => x"00000000",	--0034
0014 => x"00000000",	--0038
0015 => x"00000000",	--003C
0016 => x"00000000",	--0040
0017 => x"00000000",	--0044
0018 => x"00000000",	--0048
0019 => x"00000000",	--004C
0020 => x"00000000",	--0050
0021 => x"00000000",	--0054
0022 => x"00000000",	--0058
0023 => x"00000000",	--005C
0024 => x"00000000",	--0060
0025 => x"00000000",	--0064
0026 => x"00000000",	--0068
0027 => x"00000000",	--006C
0028 => x"00000000",	--0070
0029 => x"00000000",	--0074
0030 => x"00000000",	--0078
0031 => x"00000000",	--007C
0032 => x"00000000",	--0080
0033 => x"00000000",	--0084
0034 => x"00000000",	--0088
0035 => x"00000000",	--008C
0036 => x"00000000",	--0090
0037 => x"00000000",	--0094
0038 => x"00000000",	--0098
0039 => x"00000000",	--009C
0040 => x"00000000",	--00A0
0041 => x"00000000",	--00A4
0042 => x"60020101",	--00A8
0043 => x"60040001",	--00AC
0044 => x"60010020",	--00B0
0045 => x"80000008",	--00B4
0046 => x"64880040",	--00B8
0047 => x"64820140",	--00BC
0048 => x"80000010",	--00C0
0049 => x"64820140",	--00C4
0050 => x"80000010",	--00C8
0051 => x"64860140",	--00CC
0052 => x"80000077",	--00D0
0053 => x"648A0140",	--00D4
0054 => x"400000D0",	--00D8
0055 => x"800000A0",	--00DC
0056 => x"602C0000",	--00E0
0057 => x"64800040",	--00E4
0058 => x"60003040",	--00E8
0059 => x"64020140",	--00EC
0060 => x"400000D0",	--00F0
0061 => x"800000A0",	--00F4
0062 => x"602C0000",	--00F8
0063 => x"64800040",	--00FC
0064 => x"602E1100",	--0100
0065 => x"80000020",	--0104
0066 => x"80000080",	--0108
0067 => x"80000000",	--010C
0068 => x"00000918",	--0110
0069 => x"80000008",	--0114
0070 => x"640080C0",	--0118
0071 => x"80000000",	--011C
0072 => x"640080C0",	--0120
0073 => x"68010020",	--0124
0074 => x"80000003",	--0128
0075 => x"60000001",	--012C
0076 => x"64A80040",	--0130
0077 => x"64010020",	--0134
0078 => x"40000910",	--0138
0079 => x"68000021",	--013C
0080 => x"6C988000",	--0140
0081 => x"20000124",	--0144
0082 => x"60000100",	--0148
0083 => x"60000100",	--014C
0084 => x"64020140",	--0150
0085 => x"800000A0",	--0154
0086 => x"602C0000",	--0158
0087 => x"64800040",	--015C
0088 => x"80000008",	--0160
0089 => x"64800000",	--0164
0090 => x"64010000",	--0168
0091 => x"64010000",	--016C
0092 => x"640080C0",	--0170
0093 => x"640080C0",	--0174
0094 => x"68010020",	--0178
0095 => x"602C1000",	--017C
0096 => x"2000018C",	--0180
0097 => x"80000023",	--0184
0098 => x"00000190",	--0188
0099 => x"8000002E",	--018C
0100 => x"40000800",	--0190
0101 => x"80000020",	--0194
0102 => x"40000800",	--0198
0103 => x"68000021",	--019C
0104 => x"6C988000",	--01A0
0105 => x"20000178",	--01A4
0106 => x"60000100",	--01A8
0107 => x"60000100",	--01AC
0108 => x"0000081C",	--01B0
0109 => x"80000154",	--01B4
0110 => x"00000114",	--01B8
0111 => x"60010020",	--01BC
0112 => x"400000AC",	--01C0
0113 => x"400000C8",	--01C4
0114 => x"400000F0",	--01C8
0115 => x"64010020",	--01CC
0116 => x"400000C8",	--01D0
0117 => x"400000F0",	--01D4
0118 => x"64800040",	--01D8
0119 => x"64010020",	--01DC
0120 => x"400000A8",	--01E0
0121 => x"400000C8",	--01E4
0122 => x"400000F0",	--01E8
0123 => x"64800040",	--01EC
0124 => x"64010020",	--01F0
0125 => x"400000AC",	--01F4
0126 => x"400000F0",	--01F8
0127 => x"64800040",	--01FC
0128 => x"64010020",	--0200
0129 => x"400000A8",	--0204
0130 => x"400000F0",	--0208
0131 => x"64800040",	--020C
0132 => x"64010020",	--0210
0133 => x"400000AC",	--0214
0134 => x"400000C0",	--0218
0135 => x"400000F0",	--021C
0136 => x"64800040",	--0220
0137 => x"64010020",	--0224
0138 => x"400000C0",	--0228
0139 => x"400000F0",	--022C
0140 => x"64800040",	--0230
0141 => x"64010020",	--0234
0142 => x"400000A8",	--0238
0143 => x"400000C0",	--023C
0144 => x"400000F0",	--0240
0145 => x"64820140",	--0244
0146 => x"400001BC",	--0248
0147 => x"64010020",	--024C
0148 => x"800000A0",	--0250
0149 => x"602C0000",	--0254
0150 => x"64800040",	--0258
0151 => x"602C1000",	--025C
0152 => x"648C0040",	--0260
0153 => x"80000003",	--0264
0154 => x"64980040",	--0268
0155 => x"80000001",	--026C
0156 => x"64880040",	--0270
0157 => x"64010000",	--0274
0158 => x"800000A4",	--0278
0159 => x"602C0000",	--027C
0160 => x"64800040",	--0280
0161 => x"60003040",	--0284
0162 => x"64020140",	--0288
0163 => x"80000008",	--028C
0164 => x"64800000",	--0290
0165 => x"64010000",	--0294
0166 => x"64010000",	--0298
0167 => x"640080C0",	--029C
0168 => x"640080C0",	--02A0
0169 => x"68010020",	--02A4
0170 => x"40000248",	--02A8
0171 => x"68000021",	--02AC
0172 => x"6C988000",	--02B0
0173 => x"200002A4",	--02B4
0174 => x"60000100",	--02B8
0175 => x"60000100",	--02BC
0176 => x"60020100",	--02C0
0177 => x"800000A0",	--02C4
0178 => x"602C0000",	--02C8
0179 => x"800000A4",	--02CC
0180 => x"602C0000",	--02D0
0181 => x"800000A0",	--02D4
0182 => x"60002040",	--02D8
0183 => x"64000040",	--02DC
0184 => x"800000A4",	--02E0
0185 => x"60002040",	--02E4
0186 => x"64020140",	--02E8
0187 => x"8000028C",	--02EC
0188 => x"40000114",	--02F0
0189 => x"000002C4",	--02F4
0190 => x"640080C0",	--02F8
0191 => x"64010000",	--02FC
0192 => x"68010120",	--0300
0193 => x"64010000",	--0304
0194 => x"60010020",	--0308
0195 => x"40000874",	--030C
0196 => x"64800000",	--0310
0197 => x"64010000",	--0314
0198 => x"64010000",	--0318
0199 => x"640080C0",	--031C
0200 => x"640080C0",	--0320
0201 => x"68010020",	--0324
0202 => x"602C1000",	--0328
0203 => x"8000007C",	--032C
0204 => x"64980040",	--0330
0205 => x"20000348",	--0334
0206 => x"64000040",	--0338
0207 => x"400000C0",	--033C
0208 => x"60010020",	--0340
0209 => x"00000368",	--0344
0210 => x"68010020",	--0348
0211 => x"602C1000",	--034C
0212 => x"80000020",	--0350
0213 => x"64980040",	--0354
0214 => x"60000001",	--0358
0215 => x"64010020",	--035C
0216 => x"400000D8",	--0360
0217 => x"400000A8",	--0364
0218 => x"68000021",	--0368
0219 => x"6C988000",	--036C
0220 => x"20000324",	--0370
0221 => x"60000100",	--0374
0222 => x"60000100",	--0378
0223 => x"000008A0",	--037C
0224 => x"400008F0",	--0380
0225 => x"7C2A200A",	--0384
0226 => x"7C2A2020",	--0388
0227 => x"002A2A2A",	--038C
0228 => x"000002F8",	--0390
0229 => x"400008F0",	--0394
0230 => x"2A2A2A03",	--0398
0231 => x"000002F8",	--039C
0232 => x"80000020",	--03A0
0233 => x"800000A0",	--03A4
0234 => x"60002040",	--03A8
0235 => x"64000040",	--03AC
0236 => x"80000020",	--03B0
0237 => x"80000008",	--03B4
0238 => x"64800040",	--03B8
0239 => x"800000A4",	--03BC
0240 => x"60002040",	--03C0
0241 => x"64000040",	--03C4
0242 => x"80000003",	--03C8
0243 => x"40000380",	--03CC
0244 => x"400001B4",	--03D0
0245 => x"4000081C",	--03D4
0246 => x"400002EC",	--03D8
0247 => x"000003D0",	--03DC

0512 => x"80010000",	--0800
0513 => x"60002040",	--0804
0514 => x"64000040",	--0808
0515 => x"80010004",	--080C
0516 => x"602D0020",	--0810
0517 => x"20000810",	--0814
0518 => x"64020140",	--0818
0519 => x"8000000A",	--081C
0520 => x"00000800",	--0820
0521 => x"80000020",	--0824
0522 => x"00000800",	--0828
0523 => x"64800000",	--082C
0524 => x"64010000",	--0830
0525 => x"64010000",	--0834
0526 => x"640080C0",	--0838
0527 => x"640080C0",	--083C
0528 => x"68010020",	--0840
0529 => x"602C1000",	--0844
0530 => x"40000800",	--0848
0531 => x"68000021",	--084C
0532 => x"6C988000",	--0850
0533 => x"20000840",	--0854
0534 => x"60000100",	--0858
0535 => x"60000100",	--085C
0536 => x"60020100",	--0860
0537 => x"60010020",	--0864
0538 => x"60000001",	--0868
0539 => x"64010000",	--086C
0540 => x"602E1100",	--0870
0541 => x"640080C0",	--0874
0542 => x"64010000",	--0878
0543 => x"68010120",	--087C
0544 => x"64010000",	--0880
0545 => x"640080C0",	--0884
0546 => x"640080C0",	--0888
0547 => x"64010000",	--088C
0548 => x"68010120",	--0890
0549 => x"64010000",	--0894
0550 => x"68010120",	--0898
0551 => x"60020100",	--089C
0552 => x"64000040",	--08A0
0553 => x"64020140",	--08A4
0554 => x"60010020",	--08A8
0555 => x"200008B4",	--08AC
0556 => x"60010020",	--08B0
0557 => x"60020100",	--08B4
0558 => x"60140000",	--08B8
0559 => x"60020101",	--08BC
0560 => x"64010020",	--08C0
0561 => x"64010020",	--08C4
0562 => x"649C0040",	--08C8
0563 => x"200008D8",	--08CC
0564 => x"64000040",	--08D0
0565 => x"000008DC",	--08D4
0566 => x"60000040",	--08D8
0567 => x"60020100",	--08DC
0568 => x"64010020",	--08E0
0569 => x"64010020",	--08E4
0570 => x"611C0040",	--08E8
0571 => x"000008CC",	--08EC
0572 => x"68000020",	--08F0
0573 => x"602C1000",	--08F4
0574 => x"68810020",	--08F8
0575 => x"60240002",	--08FC
0576 => x"60280002",	--0900
0577 => x"60000004",	--0904
0578 => x"68008001",	--0908
0579 => x"64030100",	--090C
0580 => x"640080C0",	--0910
0581 => x"60020100",	--0914
0582 => x"640080C0",	--0918
0583 => x"64800000",	--091C
0584 => x"64010000",	--0920
0585 => x"64910020",	--0924
0586 => x"20000944",	--0928
0587 => x"68010020",	--092C
0588 => x"64010020",	--0930
0589 => x"60003040",	--0934
0590 => x"64000040",	--0938
0591 => x"60000001",	--093C
0592 => x"00000924",	--0940
0593 => x"68010120",	--0944
0594 => x"64000040",	--0948
0595 => x"000008A0",	--094C
0596 => x"80000000",	--0950
0597 => x"64010000",	--0954
0598 => x"640080C0",	--0958
0599 => x"640080C0",	--095C
0600 => x"64010020",	--0960
0601 => x"602C0000",	--0964
0602 => x"64010020",	--0968
0603 => x"60002040",	--096C
0604 => x"64000040",	--0970
0605 => x"60000002",	--0974
0606 => x"64010000",	--0978
0607 => x"60000002",	--097C
0608 => x"64010000",	--0980
0609 => x"68000021",	--0984
0610 => x"6C988000",	--0988
0611 => x"20000960",	--098C
0612 => x"60000100",	--0990
0613 => x"60000100",	--0994
0614 => x"000008A0",	--0998
0615 => x"80000000",	--099C
0616 => x"64010000",	--09A0
0617 => x"640080C0",	--09A4
0618 => x"640080C0",	--09A8
0619 => x"64010020",	--09AC
0620 => x"602C1000",	--09B0
0621 => x"64010020",	--09B4
0622 => x"60003040",	--09B8
0623 => x"64000040",	--09BC
0624 => x"60000001",	--09C0
0625 => x"64010000",	--09C4
0626 => x"60000001",	--09C8
0627 => x"64010000",	--09CC
0628 => x"68000021",	--09D0
0629 => x"6C988000",	--09D4
0630 => x"200009AC",	--09D8
0631 => x"60000100",	--09DC
0632 => x"60000100",	--09E0
0633 => x"000008A0",	--09E4
0634 => x"60020100",	--09E8
0635 => x"60280001",	--09EC
0636 => x"64010020",	--09F0
0637 => x"601C0000",	--09F4
0638 => x"20000A00",	--09F8
0639 => x"60000001",	--09FC
0640 => x"64290001",	--0A00
0641 => x"64010000",	--0A04
0642 => x"640080C0",	--0A08
0643 => x"64010000",	--0A0C
0644 => x"68010120",	--0A10
0645 => x"64010000",	--0A14
0646 => x"64010020",	--0A18
0647 => x"64010020",	--0A1C
0648 => x"649C0040",	--0A20
0649 => x"60140000",	--0A24
0650 => x"20000A5C",	--0A28
0651 => x"64850000",	--0A2C
0652 => x"64010000",	--0A30
0653 => x"640080C0",	--0A34
0654 => x"64010000",	--0A38
0655 => x"68010120",	--0A3C
0656 => x"64010000",	--0A40
0657 => x"60000001",	--0A44
0658 => x"640080C0",	--0A48
0659 => x"64010000",	--0A4C
0660 => x"68010120",	--0A50
0661 => x"64010000",	--0A54
0662 => x"00000A6C",	--0A58
0663 => x"64010000",	--0A5C
0664 => x"640080C0",	--0A60
0665 => x"64010000",	--0A64
0666 => x"68010120",	--0A68
0667 => x"60020100",	--0A6C
0668 => x"64010000",	--0A70
0669 => x"640080C0",	--0A74
0670 => x"64010000",	--0A78
0671 => x"68010120",	--0A7C
0672 => x"80000020",	--0A80
0673 => x"640080C0",	--0A84
0674 => x"80000000",	--0A88
0675 => x"640080C0",	--0A8C
0676 => x"400009EC",	--0A90
0677 => x"68000021",	--0A94
0678 => x"6C988000",	--0A98
0679 => x"20000A90",	--0A9C
0680 => x"60000100",	--0AA0
0681 => x"60000100",	--0AA4
0682 => x"640080C0",	--0AA8
0683 => x"64010000",	--0AAC
0684 => x"68010120",	--0AB0
0685 => x"64010000",	--0AB4
0686 => x"64000040",	--0AB8
0687 => x"64030100",	--0ABC
0688 => x"64010000",	--0AC0
0689 => x"640080C0",	--0AC4
0690 => x"64010000",	--0AC8
0691 => x"68010120",	--0ACC
0692 => x"80000020",	--0AD0
0693 => x"640080C0",	--0AD4
0694 => x"80000000",	--0AD8
0695 => x"640080C0",	--0ADC
0696 => x"400009EC",	--0AE0
0697 => x"68000021",	--0AE4
0698 => x"6C988000",	--0AE8
0699 => x"20000AE0",	--0AEC
0700 => x"60000100",	--0AF0
0701 => x"60000100",	--0AF4
0702 => x"640080C0",	--0AF8
0703 => x"64010000",	--0AFC
0704 => x"68010120",	--0B00
0705 => x"64010000",	--0B04
0706 => x"64000040",	--0B08
0707 => x"64020140",	--0B0C
0708 => x"0000000A",	--0B10
0709 => x"00000000",	--0B14
0710 => x"00000000",	--0B18
0711 => x"00000000",	--0B1C
0712 => x"00000000",	--0B20
0713 => x"00000000",	--0B24
0714 => x"00000000",	--0B28
0715 => x"00000000",	--0B2C
0716 => x"00000000",	--0B30
0717 => x"00000000",	--0B34
0718 => x"00000000",	--0B38
0719 => x"00000000",	--0B3C
0720 => x"00000000",	--0B40
0721 => x"00000000",	--0B44
0722 => x"00000000",	--0B48
0723 => x"00000000",	--0B4C
0724 => x"00000000",	--0B50
0725 => x"00000000",	--0B54
0726 => x"00000000",	--0B58
0727 => x"00000000",	--0B5C
0728 => x"00000000",	--0B60
0729 => x"00000000",	--0B64
0730 => x"00000000",	--0B68
0731 => x"80000B14",	--0B6C
0732 => x"602C0000",	--0B70
0733 => x"60040001",	--0B74
0734 => x"60010020",	--0B78
0735 => x"80000B14",	--0B7C
0736 => x"60002040",	--0B80
0737 => x"64000040",	--0B84
0738 => x"60003040",	--0B88
0739 => x"64020140",	--0B8C
0740 => x"80000009",	--0B90
0741 => x"64010020",	--0B94
0742 => x"649C0040",	--0B98
0743 => x"20000BA8",	--0B9C
0744 => x"80000007",	--0BA0
0745 => x"64800040",	--0BA4
0746 => x"80000030",	--0BA8
0747 => x"64820140",	--0BAC
0748 => x"80000B6C",	--0BB0
0749 => x"80000B14",	--0BB4
0750 => x"60002040",	--0BB8
0751 => x"64020140",	--0BBC
0752 => x"80000B10",	--0BC0
0753 => x"602C0000",	--0BC4
0754 => x"40000A70",	--0BC8
0755 => x"64010000",	--0BCC
0756 => x"40000B90",	--0BD0
0757 => x"40000B6C",	--0BD4
0758 => x"80000000",	--0BD8
0759 => x"60020100",	--0BDC
0760 => x"40000BC0",	--0BE0
0761 => x"64010020",	--0BE4
0762 => x"64010020",	--0BE8
0763 => x"648C0040",	--0BEC
0764 => x"60180000",	--0BF0
0765 => x"20000BE0",	--0BF4
0766 => x"60020100",	--0BF8
0767 => x"400008A0",	--0BFC
0768 => x"80000B14",	--0C00
0769 => x"602C0000",	--0C04
0770 => x"80000B6C",	--0C08
0771 => x"64010020",	--0C0C
0772 => x"64860140",	--0C10
0773 => x"8000000A",	--0C14
0774 => x"80000B10",	--0C18
0775 => x"60002040",	--0C1C
0776 => x"64020140",	--0C20
0777 => x"80000010",	--0C24
0778 => x"80000B10",	--0C28
0779 => x"60002040",	--0C2C
0780 => x"64020140",	--0C30

others => x"00000000"
);

begin

    a_addr_word <= a_addr(addr_bits-1 downto 2);
    b_addr_word <= b_addr(addr_bits-1 downto 2);

    process (clk, rst, a_addr_word, a_we, b_addr_word, b_we) begin
	if rising_edge(clk) then
	    if rst = '1' then
		a_dout <= (others => '0');
		b_dout <= (others => '0');
	    else
		-- Port A

		if (a_we = '1') then
		    ram(to_integer(unsigned(a_addr_word))) <= a_din;
		end if;

		a_dout <= ram(to_integer(unsigned(a_addr_word)));

		-- Port B

		if b_we(0) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(7 downto 0) <= b_din(7 downto 0);
		end if;

		if b_we(1) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(15 downto 8) <= b_din(15 downto 8);
		end if;

		if b_we(2) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(23 downto 16) <= b_din(23 downto 16);
		end if;

		if b_we(3) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(31 downto 24) <= b_din(31 downto 24);
		end if;

		b_dout <= ram(to_integer(unsigned(b_addr_word)));

	    end if;
	end if;
    end process;

end;
