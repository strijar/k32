../ghdl/ram.vhd