--
--  Copyright 2015 Oleg Belousov <belousov.oleg@gmail.com>,
--
--  All rights reserved.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--    1. Redistributions of source code must retain the above copyright notice,
--       this list of conditions and the following disclaimer.
-- 
--    2. Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.k32_pkg.all;

entity ram is
    generic (
	addr_bits	: integer := 5;
	data_bits	: integer := 16
    );
    port (
	clk	: in std_logic;
	rst	: in std_logic;

	a_addr	: in std_logic_vector(addr_bits-1 downto 0);
	a_din	: in std_logic_vector(data_bits-1 downto 0);
	a_dout	: out std_logic_vector(data_bits-1 downto 0);
        a_we	: in std_logic;

	b_en	: in std_logic;
	b_addr	: in std_logic_vector(addr_bits-1 downto 0);
	b_din	: in std_logic_vector(data_bits-1 downto 0);
	b_dout	: out std_logic_vector(data_bits-1 downto 0);
        b_we	: in std_logic_vector(3 downto 0)
    );
end ram;

architecture rtl of ram is

type ram_type is array(natural range 0 to (2**(addr_bits))-1) of std_logic_vector(data_bits-1 downto 0);

signal a_addr_word	: std_logic_vector(addr_bits-1 downto 2) := (others => '0');
signal b_addr_word	: std_logic_vector(addr_bits-1 downto 2) := (others => '0');

signal ram : ram_type :=
(
0000 => x"00000514",	--0000
0001 => x"000009E8",	--0004

0008 => x"00000000",	--0020
0009 => x"00000000",	--0024
0010 => x"00000000",	--0028
0011 => x"00000000",	--002C
0012 => x"00000000",	--0030
0013 => x"00000000",	--0034
0014 => x"00000000",	--0038
0015 => x"00000000",	--003C
0016 => x"00000000",	--0040
0017 => x"00000000",	--0044
0018 => x"00000000",	--0048
0019 => x"00000000",	--004C
0020 => x"00000000",	--0050
0021 => x"00000000",	--0054
0022 => x"00000000",	--0058
0023 => x"00000000",	--005C
0024 => x"00000000",	--0060
0025 => x"00000000",	--0064
0026 => x"00000000",	--0068
0027 => x"00000000",	--006C
0028 => x"00000000",	--0070
0029 => x"00000000",	--0074
0030 => x"00000000",	--0078
0031 => x"00000000",	--007C
0032 => x"00000000",	--0080
0033 => x"00000000",	--0084
0034 => x"00000000",	--0088
0035 => x"00000000",	--008C
0036 => x"00000000",	--0090
0037 => x"00000000",	--0094
0038 => x"00000000",	--0098
0039 => x"00000000",	--009C
0040 => x"00000000",	--00A0
0041 => x"00000000",	--00A4
0042 => x"00000000",	--00A8
0043 => x"00000000",	--00AC
0044 => x"00000000",	--00B0
0045 => x"00000000",	--00B4
0046 => x"00000000",	--00B8
0047 => x"00000000",	--00BC
0048 => x"00000000",	--00C0
0049 => x"00000000",	--00C4
0050 => x"00000000",	--00C8
0051 => x"00000000",	--00CC
0052 => x"00000000",	--00D0
0053 => x"00000000",	--00D4
0054 => x"00000000",	--00D8
0055 => x"00000000",	--00DC
0056 => x"00000000",	--00E0
0057 => x"00000000",	--00E4
0058 => x"00000000",	--00E8
0059 => x"00000000",	--00EC
0060 => x"00000000",	--00F0
0061 => x"00000000",	--00F4
0062 => x"00000000",	--00F8
0063 => x"00000000",	--00FC
0064 => x"00000000",	--0100
0065 => x"00000000",	--0104
0066 => x"00000000",	--0108
0067 => x"00000000",	--010C
0068 => x"00000000",	--0110
0069 => x"00000000",	--0114
0070 => x"00000000",	--0118
0071 => x"00000000",	--011C
0072 => x"00000000",	--0120
0073 => x"00000000",	--0124
0074 => x"00000000",	--0128
0075 => x"00000000",	--012C
0076 => x"00000000",	--0130
0077 => x"00000000",	--0134
0078 => x"00000000",	--0138
0079 => x"00000000",	--013C
0080 => x"00000000",	--0140
0081 => x"00000000",	--0144
0082 => x"00000000",	--0148
0083 => x"00000000",	--014C
0084 => x"00000000",	--0150
0085 => x"00000000",	--0154
0086 => x"00000000",	--0158
0087 => x"00000000",	--015C
0088 => x"00000000",	--0160
0089 => x"00000000",	--0164
0090 => x"00000000",	--0168
0091 => x"00000000",	--016C
0092 => x"00000000",	--0170
0093 => x"00000000",	--0174
0094 => x"00000000",	--0178
0095 => x"00000000",	--017C
0096 => x"00000000",	--0180
0097 => x"00000000",	--0184
0098 => x"00000000",	--0188
0099 => x"00000000",	--018C
0100 => x"00000000",	--0190
0101 => x"00000000",	--0194
0102 => x"00000000",	--0198
0103 => x"00000000",	--019C
0104 => x"00000000",	--01A0
0105 => x"00000000",	--01A4
0106 => x"00000000",	--01A8
0107 => x"00000000",	--01AC
0108 => x"00000000",	--01B0
0109 => x"00000000",	--01B4
0110 => x"00000000",	--01B8
0111 => x"00000000",	--01BC
0112 => x"00000000",	--01C0
0113 => x"00000000",	--01C4
0114 => x"00000000",	--01C8
0115 => x"00000000",	--01CC
0116 => x"00000000",	--01D0
0117 => x"00000000",	--01D4
0118 => x"00000000",	--01D8
0119 => x"00000000",	--01DC
0120 => x"00000000",	--01E0
0121 => x"00000000",	--01E4
0122 => x"00000000",	--01E8
0123 => x"00000000",	--01EC
0124 => x"00000000",	--01F0
0125 => x"00000000",	--01F4
0126 => x"00000000",	--01F8
0127 => x"00000000",	--01FC
0128 => x"00000000",	--0200
0129 => x"00000000",	--0204
0130 => x"00000000",	--0208
0131 => x"00000000",	--020C
0132 => x"00000000",	--0210
0133 => x"00000000",	--0214
0134 => x"00000000",	--0218
0135 => x"00000000",	--021C
0136 => x"00000000",	--0220
0137 => x"00000000",	--0224
0138 => x"60080201",	--0228
0139 => x"60100001",	--022C
0140 => x"60040020",	--0230
0141 => x"80000010",	--0234
0142 => x"65200040",	--0238
0143 => x"65080240",	--023C
0144 => x"80000020",	--0240
0145 => x"65080240",	--0244
0146 => x"80000020",	--0248
0147 => x"65180240",	--024C
0148 => x"800001EF",	--0250
0149 => x"65280240",	--0254
0150 => x"40000250",	--0258
0151 => x"80000220",	--025C
0152 => x"60B00000",	--0260
0153 => x"65000040",	--0264
0154 => x"60018040",	--0268
0155 => x"64080240",	--026C
0156 => x"40000250",	--0270
0157 => x"80000220",	--0274
0158 => x"60B00000",	--0278
0159 => x"65000040",	--027C
0160 => x"60B88200",	--0280
0161 => x"80000020",	--0284
0162 => x"80000200",	--0288
0163 => x"80000000",	--028C
0164 => x"00000918",	--0290
0165 => x"80000010",	--0294
0166 => x"64020140",	--0298
0167 => x"80000000",	--029C
0168 => x"64020140",	--02A0
0169 => x"68040020",	--02A4
0170 => x"80000004",	--02A8
0171 => x"60000001",	--02AC
0172 => x"65A00040",	--02B0
0173 => x"64040020",	--02B4
0174 => x"40000910",	--02B8
0175 => x"68000021",	--02BC
0176 => x"6D620000",	--02C0
0177 => x"200002A4",	--02C4
0178 => x"60000200",	--02C8
0179 => x"60000200",	--02CC
0180 => x"64080240",	--02D0
0181 => x"80000220",	--02D4
0182 => x"60B00000",	--02D8
0183 => x"65000040",	--02DC
0184 => x"80000010",	--02E0
0185 => x"65000000",	--02E4
0186 => x"64040000",	--02E8
0187 => x"64040000",	--02EC
0188 => x"64020140",	--02F0
0189 => x"64020140",	--02F4
0190 => x"68040020",	--02F8
0191 => x"60B08000",	--02FC
0192 => x"2000030C",	--0300
0193 => x"80000023",	--0304
0194 => x"00000310",	--0308
0195 => x"8000002E",	--030C
0196 => x"40000800",	--0310
0197 => x"80000020",	--0314
0198 => x"40000800",	--0318
0199 => x"68000021",	--031C
0200 => x"6D620000",	--0320
0201 => x"200002F8",	--0324
0202 => x"60000200",	--0328
0203 => x"60000200",	--032C
0204 => x"0000081C",	--0330
0205 => x"800002D4",	--0334
0206 => x"00000294",	--0338
0207 => x"60040020",	--033C
0208 => x"4000022C",	--0340
0209 => x"40000248",	--0344
0210 => x"40000270",	--0348
0211 => x"64040020",	--034C
0212 => x"40000248",	--0350
0213 => x"40000270",	--0354
0214 => x"65000040",	--0358
0215 => x"64040020",	--035C
0216 => x"40000228",	--0360
0217 => x"40000248",	--0364
0218 => x"40000270",	--0368
0219 => x"65000040",	--036C
0220 => x"64040020",	--0370
0221 => x"4000022C",	--0374
0222 => x"40000270",	--0378
0223 => x"65000040",	--037C
0224 => x"64040020",	--0380
0225 => x"40000228",	--0384
0226 => x"40000270",	--0388
0227 => x"65000040",	--038C
0228 => x"64040020",	--0390
0229 => x"4000022C",	--0394
0230 => x"40000240",	--0398
0231 => x"40000270",	--039C
0232 => x"65000040",	--03A0
0233 => x"64040020",	--03A4
0234 => x"40000240",	--03A8
0235 => x"40000270",	--03AC
0236 => x"65000040",	--03B0
0237 => x"64040020",	--03B4
0238 => x"40000228",	--03B8
0239 => x"40000240",	--03BC
0240 => x"40000270",	--03C0
0241 => x"65080240",	--03C4
0242 => x"4000033C",	--03C8
0243 => x"64040020",	--03CC
0244 => x"80000220",	--03D0
0245 => x"60B00000",	--03D4
0246 => x"65000040",	--03D8
0247 => x"60B08000",	--03DC
0248 => x"65300040",	--03E0
0249 => x"80000003",	--03E4
0250 => x"65600040",	--03E8
0251 => x"80000001",	--03EC
0252 => x"65200040",	--03F0
0253 => x"64040000",	--03F4
0254 => x"80000224",	--03F8
0255 => x"60B00000",	--03FC
0256 => x"65000040",	--0400
0257 => x"60018040",	--0404
0258 => x"64080240",	--0408
0259 => x"80000010",	--040C
0260 => x"65000000",	--0410
0261 => x"64040000",	--0414
0262 => x"64040000",	--0418
0263 => x"64020140",	--041C
0264 => x"64020140",	--0420
0265 => x"68040020",	--0424
0266 => x"400003C8",	--0428
0267 => x"68000021",	--042C
0268 => x"6D620000",	--0430
0269 => x"20000424",	--0434
0270 => x"60000200",	--0438
0271 => x"60000200",	--043C
0272 => x"60080200",	--0440
0273 => x"80000220",	--0444
0274 => x"60B00000",	--0448
0275 => x"80000224",	--044C
0276 => x"60B00000",	--0450
0277 => x"80000220",	--0454
0278 => x"60010040",	--0458
0279 => x"64000040",	--045C
0280 => x"80000224",	--0460
0281 => x"60010040",	--0464
0282 => x"64080240",	--0468
0283 => x"8000040C",	--046C
0284 => x"40000294",	--0470
0285 => x"00000444",	--0474
0286 => x"64020140",	--0478
0287 => x"64040000",	--047C
0288 => x"68040220",	--0480
0289 => x"64040000",	--0484
0290 => x"60040020",	--0488
0291 => x"40000874",	--048C
0292 => x"65000000",	--0490
0293 => x"64040000",	--0494
0294 => x"64040000",	--0498
0295 => x"64020140",	--049C
0296 => x"64020140",	--04A0
0297 => x"68040020",	--04A4
0298 => x"60B08000",	--04A8
0299 => x"8000007C",	--04AC
0300 => x"65600040",	--04B0
0301 => x"200004C8",	--04B4
0302 => x"64000040",	--04B8
0303 => x"40000240",	--04BC
0304 => x"60040020",	--04C0
0305 => x"000004E8",	--04C4
0306 => x"68040020",	--04C8
0307 => x"60B08000",	--04CC
0308 => x"80000020",	--04D0
0309 => x"65600040",	--04D4
0310 => x"60000001",	--04D8
0311 => x"64040020",	--04DC
0312 => x"40000258",	--04E0
0313 => x"40000228",	--04E4
0314 => x"68000021",	--04E8
0315 => x"6D620000",	--04EC
0316 => x"200004A4",	--04F0
0317 => x"60000200",	--04F4
0318 => x"60000200",	--04F8
0319 => x"000008A0",	--04FC
0320 => x"400008F0",	--0500
0321 => x"7C2A200A",	--0504
0322 => x"7C2A2020",	--0508
0323 => x"002A2A2A",	--050C
0324 => x"00000478",	--0510
0325 => x"80000020",	--0514
0326 => x"80000220",	--0518
0327 => x"60010040",	--051C
0328 => x"64000040",	--0520
0329 => x"80000020",	--0524
0330 => x"80000010",	--0528
0331 => x"65000040",	--052C
0332 => x"80000224",	--0530
0333 => x"60010040",	--0534
0334 => x"64000040",	--0538
0335 => x"80000000",	--053C
0336 => x"40000500",	--0540
0337 => x"40000334",	--0544
0338 => x"4000081C",	--0548
0339 => x"4000046C",	--054C
0340 => x"00000544",	--0550

0512 => x"80010000",	--0800
0513 => x"60010040",	--0804
0514 => x"64000040",	--0808
0515 => x"80010004",	--080C
0516 => x"60B40020",	--0810
0517 => x"20000810",	--0814
0518 => x"64080240",	--0818
0519 => x"8000000A",	--081C
0520 => x"00000800",	--0820
0521 => x"80000020",	--0824
0522 => x"00000800",	--0828
0523 => x"65000000",	--082C
0524 => x"64040000",	--0830
0525 => x"64040000",	--0834
0526 => x"64020140",	--0838
0527 => x"64020140",	--083C
0528 => x"68040020",	--0840
0529 => x"60B08000",	--0844
0530 => x"40000800",	--0848
0531 => x"68000021",	--084C
0532 => x"6D620000",	--0850
0533 => x"20000840",	--0854
0534 => x"60000200",	--0858
0535 => x"60000200",	--085C
0536 => x"60080200",	--0860
0537 => x"60040020",	--0864
0538 => x"60000001",	--0868
0539 => x"64040000",	--086C
0540 => x"60B88200",	--0870
0541 => x"64020140",	--0874
0542 => x"64040000",	--0878
0543 => x"68040220",	--087C
0544 => x"64040000",	--0880
0545 => x"64020140",	--0884
0546 => x"64020140",	--0888
0547 => x"64040000",	--088C
0548 => x"68040220",	--0890
0549 => x"64040000",	--0894
0550 => x"68040220",	--0898
0551 => x"60080200",	--089C
0552 => x"64000040",	--08A0
0553 => x"64080240",	--08A4
0554 => x"60040020",	--08A8
0555 => x"200008B4",	--08AC
0556 => x"60040020",	--08B0
0557 => x"60080200",	--08B4
0558 => x"60500000",	--08B8
0559 => x"60080201",	--08BC
0560 => x"64040020",	--08C0
0561 => x"64040020",	--08C4
0562 => x"65700040",	--08C8
0563 => x"200008D8",	--08CC
0564 => x"64000040",	--08D0
0565 => x"000008DC",	--08D4
0566 => x"60000040",	--08D8
0567 => x"60080200",	--08DC
0568 => x"64040020",	--08E0
0569 => x"64040020",	--08E4
0570 => x"62700040",	--08E8
0571 => x"000008CC",	--08EC
0572 => x"68000020",	--08F0
0573 => x"60B08000",	--08F4
0574 => x"69040020",	--08F8
0575 => x"60900002",	--08FC
0576 => x"60A00002",	--0900
0577 => x"60000004",	--0904
0578 => x"68020001",	--0908
0579 => x"640C0200",	--090C
0580 => x"64020140",	--0910
0581 => x"60080200",	--0914
0582 => x"64020140",	--0918
0583 => x"65000000",	--091C
0584 => x"64040000",	--0920
0585 => x"65440020",	--0924
0586 => x"20000944",	--0928
0587 => x"68040020",	--092C
0588 => x"64040020",	--0930
0589 => x"60018040",	--0934
0590 => x"64000040",	--0938
0591 => x"60000001",	--093C
0592 => x"00000924",	--0940
0593 => x"68040220",	--0944
0594 => x"64000040",	--0948
0595 => x"000008A0",	--094C
0596 => x"80000000",	--0950
0597 => x"64040000",	--0954
0598 => x"64020140",	--0958
0599 => x"64020140",	--095C
0600 => x"64040020",	--0960
0601 => x"60B00000",	--0964
0602 => x"64040020",	--0968
0603 => x"60010040",	--096C
0604 => x"64000040",	--0970
0605 => x"60000002",	--0974
0606 => x"64040000",	--0978
0607 => x"60000002",	--097C
0608 => x"64040000",	--0980
0609 => x"68000021",	--0984
0610 => x"6D620000",	--0988
0611 => x"20000960",	--098C
0612 => x"60000200",	--0990
0613 => x"60000200",	--0994
0614 => x"000008A0",	--0998
0615 => x"80000000",	--099C
0616 => x"64040000",	--09A0
0617 => x"64020140",	--09A4
0618 => x"64020140",	--09A8
0619 => x"64040020",	--09AC
0620 => x"60B08000",	--09B0
0621 => x"64040020",	--09B4
0622 => x"60018040",	--09B8
0623 => x"64000040",	--09BC
0624 => x"60000001",	--09C0
0625 => x"64040000",	--09C4
0626 => x"60000001",	--09C8
0627 => x"64040000",	--09CC
0628 => x"68000021",	--09D0
0629 => x"6D620000",	--09D4
0630 => x"200009AC",	--09D8
0631 => x"60000200",	--09DC
0632 => x"60000200",	--09E0
0633 => x"000008A0",	--09E4
0634 => x"60080200",	--09E8
0635 => x"60A00001",	--09EC
0636 => x"64040020",	--09F0
0637 => x"60700000",	--09F4
0638 => x"20000A00",	--09F8
0639 => x"60000001",	--09FC
0640 => x"64A40001",	--0A00
0641 => x"64040000",	--0A04
0642 => x"64020140",	--0A08
0643 => x"64040000",	--0A0C
0644 => x"68040220",	--0A10
0645 => x"64040000",	--0A14
0646 => x"64040020",	--0A18
0647 => x"64040020",	--0A1C
0648 => x"65700040",	--0A20
0649 => x"60500000",	--0A24
0650 => x"20000A5C",	--0A28
0651 => x"65140000",	--0A2C
0652 => x"64040000",	--0A30
0653 => x"64020140",	--0A34
0654 => x"64040000",	--0A38
0655 => x"68040220",	--0A3C
0656 => x"64040000",	--0A40
0657 => x"60000001",	--0A44
0658 => x"64020140",	--0A48
0659 => x"64040000",	--0A4C
0660 => x"68040220",	--0A50
0661 => x"64040000",	--0A54
0662 => x"00000A6C",	--0A58
0663 => x"64040000",	--0A5C
0664 => x"64020140",	--0A60
0665 => x"64040000",	--0A64
0666 => x"68040220",	--0A68
0667 => x"60080200",	--0A6C
0668 => x"64040000",	--0A70
0669 => x"64020140",	--0A74
0670 => x"64040000",	--0A78
0671 => x"68040220",	--0A7C
0672 => x"80000020",	--0A80
0673 => x"64020140",	--0A84
0674 => x"80000000",	--0A88
0675 => x"64020140",	--0A8C
0676 => x"400009EC",	--0A90
0677 => x"68000021",	--0A94
0678 => x"6D620000",	--0A98
0679 => x"20000A90",	--0A9C
0680 => x"60000200",	--0AA0
0681 => x"60000200",	--0AA4
0682 => x"64020140",	--0AA8
0683 => x"64040000",	--0AAC
0684 => x"68040220",	--0AB0
0685 => x"64040000",	--0AB4
0686 => x"64000040",	--0AB8
0687 => x"640C0200",	--0ABC
0688 => x"64040000",	--0AC0
0689 => x"64020140",	--0AC4
0690 => x"64040000",	--0AC8
0691 => x"68040220",	--0ACC
0692 => x"80000020",	--0AD0
0693 => x"64020140",	--0AD4
0694 => x"80000000",	--0AD8
0695 => x"64020140",	--0ADC
0696 => x"400009EC",	--0AE0
0697 => x"68000021",	--0AE4
0698 => x"6D620000",	--0AE8
0699 => x"20000AE0",	--0AEC
0700 => x"60000200",	--0AF0
0701 => x"60000200",	--0AF4
0702 => x"64020140",	--0AF8
0703 => x"64040000",	--0AFC
0704 => x"68040220",	--0B00
0705 => x"64040000",	--0B04
0706 => x"64000040",	--0B08
0707 => x"64080240",	--0B0C
0708 => x"00000000",	--0B10
0709 => x"00000000",	--0B14
0710 => x"00000000",	--0B18
0711 => x"00000000",	--0B1C
0712 => x"00000000",	--0B20
0713 => x"00000000",	--0B24
0714 => x"00000000",	--0B28
0715 => x"00000000",	--0B2C
0716 => x"00000000",	--0B30
0717 => x"00000000",	--0B34
0718 => x"00000000",	--0B38
0719 => x"00000000",	--0B3C
0720 => x"00000000",	--0B40
0721 => x"00000000",	--0B44
0722 => x"00000000",	--0B48
0723 => x"00000000",	--0B4C
0724 => x"00000000",	--0B50
0725 => x"00000000",	--0B54
0726 => x"00000000",	--0B58
0727 => x"00000000",	--0B5C
0728 => x"00000000",	--0B60
0729 => x"00000000",	--0B64
0730 => x"00000000",	--0B68
0731 => x"80000B14",	--0B6C
0732 => x"60B00000",	--0B70
0733 => x"60100001",	--0B74
0734 => x"60040020",	--0B78
0735 => x"80000B14",	--0B7C
0736 => x"60010040",	--0B80
0737 => x"64000040",	--0B84
0738 => x"60018040",	--0B88
0739 => x"64080240",	--0B8C
0740 => x"80000009",	--0B90
0741 => x"64040020",	--0B94
0742 => x"65700040",	--0B98
0743 => x"20000BA8",	--0B9C
0744 => x"80000007",	--0BA0
0745 => x"65000040",	--0BA4
0746 => x"80000030",	--0BA8
0747 => x"65080240",	--0BAC
0748 => x"80000B6C",	--0BB0
0749 => x"80000B14",	--0BB4
0750 => x"60010040",	--0BB8
0751 => x"64080240",	--0BBC
0752 => x"80000B10",	--0BC0
0753 => x"60B00000",	--0BC4
0754 => x"40000A70",	--0BC8
0755 => x"64040000",	--0BCC
0756 => x"40000B90",	--0BD0
0757 => x"40000B6C",	--0BD4
0758 => x"80000000",	--0BD8
0759 => x"60080200",	--0BDC
0760 => x"40000BC0",	--0BE0
0761 => x"64040020",	--0BE4
0762 => x"64040020",	--0BE8
0763 => x"65300040",	--0BEC
0764 => x"60600000",	--0BF0
0765 => x"20000BE0",	--0BF4
0766 => x"60080200",	--0BF8
0767 => x"400008A0",	--0BFC
0768 => x"80000B14",	--0C00
0769 => x"60B00000",	--0C04
0770 => x"80000B6C",	--0C08
0771 => x"64040020",	--0C0C
0772 => x"65180240",	--0C10
0773 => x"8000000A",	--0C14
0774 => x"80000B10",	--0C18
0775 => x"60010040",	--0C1C
0776 => x"64080240",	--0C20
0777 => x"80000010",	--0C24
0778 => x"80000B10",	--0C28
0779 => x"60010040",	--0C2C
0780 => x"64080240",	--0C30
0781 => x"00000000",	--0C34
0782 => x"00000000",	--0C38
0783 => x"00000000",	--0C3C
0784 => x"00000000",	--0C40
0785 => x"00000000",	--0C44
0786 => x"00000000",	--0C48
0787 => x"00000000",	--0C4C
0788 => x"00000000",	--0C50
0789 => x"80000C54",	--0C54
0790 => x"80000C34",	--0C58
0791 => x"60010040",	--0C5C
0792 => x"64000040",	--0C60
0793 => x"78040020",	--0C64
0794 => x"60040020",	--0C68
0795 => x"60040020",	--0C6C
0796 => x"60740020",	--0C70
0797 => x"40000BB0",	--0C74
0798 => x"8000003E",	--0C78
0799 => x"40000B6C",	--0C7C
0800 => x"40000BE0",	--0C80
0801 => x"8000003C",	--0C84
0802 => x"40000B6C",	--0C88
0803 => x"40000BFC",	--0C8C
0804 => x"4000082C",	--0C90
0805 => x"40000824",	--0C94
0806 => x"400008A8",	--0C98
0807 => x"20000D48",	--0C9C
0808 => x"64020140",	--0CA0
0809 => x"80000000",	--0CA4
0810 => x"64020140",	--0CA8
0811 => x"64040000",	--0CAC
0812 => x"80000C34",	--0CB0
0813 => x"60B00000",	--0CB4
0814 => x"60100004",	--0CB8
0815 => x"60040020",	--0CBC
0816 => x"80000C34",	--0CC0
0817 => x"60010040",	--0CC4
0818 => x"64000040",	--0CC8
0819 => x"60010040",	--0CCC
0820 => x"64000040",	--0CD0
0821 => x"68000021",	--0CD4
0822 => x"6D620000",	--0CD8
0823 => x"20000CAC",	--0CDC
0824 => x"60000200",	--0CE0
0825 => x"60000200",	--0CE4
0826 => x"64020140",	--0CE8
0827 => x"80000000",	--0CEC
0828 => x"64020140",	--0CF0
0829 => x"80000C34",	--0CF4
0830 => x"60B00000",	--0CF8
0831 => x"60040020",	--0CFC
0832 => x"60000004",	--0D00
0833 => x"80000C34",	--0D04
0834 => x"60010040",	--0D08
0835 => x"64000040",	--0D0C
0836 => x"60B00000",	--0D10
0837 => x"60040020",	--0D14
0838 => x"60740020",	--0D18
0839 => x"40000BB0",	--0D1C
0840 => x"40000BE0",	--0D20
0841 => x"40000BFC",	--0D24
0842 => x"4000082C",	--0D28
0843 => x"40000824",	--0D2C
0844 => x"68000021",	--0D30
0845 => x"6D620000",	--0D34
0846 => x"20000CF4",	--0D38
0847 => x"60000200",	--0D3C
0848 => x"60000200",	--0D40
0849 => x"00000D4C",	--0D44
0850 => x"64000040",	--0D48
0851 => x"60080200",	--0D4C

others => x"00000000"
);

begin

    a_addr_word <= a_addr(addr_bits-1 downto 2);
    b_addr_word <= b_addr(addr_bits-1 downto 2);

    process (clk, rst, a_addr_word, a_we, b_addr_word, b_we) begin
	if rising_edge(clk) then
	    if rst = '1' then
		a_dout <= (others => '0');
		b_dout <= (others => '0');
	    else
		-- Port A

		if (a_we = '1') then
		    ram(to_integer(unsigned(a_addr_word))) <= a_din;
		end if;

		a_dout <= ram(to_integer(unsigned(a_addr_word)));

		-- Port B

		if b_we(0) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(7 downto 0) <= b_din(7 downto 0);
		end if;

		if b_we(1) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(15 downto 8) <= b_din(15 downto 8);
		end if;

		if b_we(2) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(23 downto 16) <= b_din(23 downto 16);
		end if;

		if b_we(3) = '1' then
		    ram(to_integer(unsigned(b_addr_word)))(31 downto 24) <= b_din(31 downto 24);
		end if;

		b_dout <= ram(to_integer(unsigned(b_addr_word)));

	    end if;
	end if;
    end process;

end;
